hiii i am iron man
